library IEEE;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity Processador_7Instrucoes is
    generic(
        WIDTH: integer := 16;
        ADDR_MSIZE: integer := 4
    );
    port (

  ) ;
end Processador_7Instrucoes;