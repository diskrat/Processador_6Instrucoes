library verilog;
use verilog.vl_types.all;
entity Processador_7Instrucoes_vlg_vec_tst is
end Processador_7Instrucoes_vlg_vec_tst;
